/*
 * Bundles up bit-encoding, bit-stuffing and nrzi
 */

// Includes
`include "nrzi.sv"
`include "stuffer.sv"
`include "crcEncoding.sv"


